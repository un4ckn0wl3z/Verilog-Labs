// Hello World Module
module hello_world ();
    // Display the message in the console on a new line with a TAB
    initial begin
        $display("\n\t Hello World! \n");
    end
endmodule